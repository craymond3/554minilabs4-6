module ab_mem_tb();

endmodule